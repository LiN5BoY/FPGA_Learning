`timescale 1ns/1ns //时间尺度、精度单位定义，决定“#（不可被综合，但在可
//综合代码中也可以写，只是会在仿真时表达效果，而综合
//时会自动被综合器优化掉）”后面的数字表示的时间尺度和
//精度，具体表达含义为:“时间尺度/时间精度”。为了以后
//编写方便我们将该句放在所有“.v”文件的开头，后面的代
//码示例将不再显示该句

module tb_mux2_1();//testbench的格式和待测试RTL模块的格式相同
//也是以“module”开始以“endmodule”结束，所有的代码都要
//在它们中间编写。不同的是在testbench中端口列表为空
//因为testbench不对外进行信号的输入输出，只是自己产生
//激励信号提供给内部实例化待测RTL模块使用，所以端口列表
//中没有内容，只是列出“()”，当然可以将“()”省略，括号
//后有个“;”不要忘记

//要在initial块和always块中被赋值的变量一定要是reg型
//在testbench中待测试RTL模块的输入永远是reg型变量
reg in1;
reg in2;
reg sel;

//输出信号，我们直接观察，也不用在任何地方进行赋值
//所以是wire型变量（在testbench中待测试RTL模块的输出永远是wire型变量）
wire out;

//initial语句是可以被综合的，一般只在testbench中表达而不在RTL代码中表达
//initial块中的语句上电后只执行一次，主要用于初始化仿真中要输入的信号
//初始化值在没有特殊要求的情况下给0或1都可以。如果不赋初值，仿真时信号
//会显示为不定态（ModelSim中的波形显示红色）
initial
begin //在仿真中begin...end块中的内容都是顺序执行的，
//在没有延时的情况下几乎没有差别，看上去是同时执行的，
//如果有延时才能表达的比较明了；
//而在rtl代码中begin...end相当于括号的作用，
//在同一个always块中给多个变量赋值的时候要加上
in1 <= 1'b0;
in2 <= 1'b0;
sel <= 1'b0;
end

//in1:产生输入随机数，模拟输入端1的输入情况
always #10 in1 <= {$random} % 2;//取模求余数，产生随机数1'b0、1'b1
//每隔10ns产生一次随机数

//in2:产生输入随机数，模拟输入端2的输入情况
always #10 in2 <= {$random} % 2;

//sel:产生输入随机数，模拟选择端的输入情况
always #10 sel <= {$random} % 2;

//下面的语句是为了在ModelSim仿真中直接打印出来信息便于观察信号变化的状态
//也可以不使用下面的语句而直接观察仿真出的波形
//------------------------------------------------------------
initial begin
$timeformat(-9, 0, "ns", 6);//设置显示的时间格式，此处表示的是(打印时间单
//位为纳秒，小数点后打印的小数位为0位，时间值
//后打印的字符串为“ns”，打印的最小数量字符为6个)

//只要监测的变量（时间、in1, in2, sel, out）发生变化，就会打印出相应的信息
$monitor("@time %t:in1=%b in2=%b sel=%b out=%b",$time,in1,in2,sel,out);
end
//------------------------------------------------------------

//待测试RTL模块的实例化，相当于将待测试模块放到测试模块中，并将输入输出对应连接上
//测试模块中产生激励信号给待测试模块的输入，以观察待测试模块的输出信号是否正确
//------------------------mux2_1_inst------------------------
mux2_1 mux2_1_inst //第一个是被实例化模块的名子，第二个是我们自己定义的在另一个
//模块中实例化后的名字。同一个模块可以在另一个模块中或不同的
//另外模块中被多次实例化，第一个名字相同，第二个名字不同
(
//前面的“in1”表示被实例化模块中的信号，后面的“in1”表示实例化该模块并要和这个
//模块的该信号相连接的信号（可以取名不同，一般取名相同，方便连接和观察）
//“.”可以理解为将这两个信号连接在一起
.in1(in1), //input in1
.in2(in2), //input in2
.sel(sel), //inputsel

.out(out) //output out
);

endmodule